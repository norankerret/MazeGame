
typedef struct packed{
	integer rowstart;
	integer colstart;
	integer width;
	integer length;	
} barrier_struct;

typedef struct packed {
	integer rowstart;
	integer colstart;
	integer width;
	integer length;
} endzone_struct;

typedef struct packed {
	integer rowstart;
	integer colstart;
	integer width;
	integer length;
} win_struct;

typedef struct packed {
	integer rowstart;
	integer colstart;
	integer width;
	integer length;
} lose_struct;

typedef struct packed {
	integer rowstart;
	integer colstart;
	integer width;
	integer length;
} confetti_struct;